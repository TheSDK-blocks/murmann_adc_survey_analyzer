*** Example netlist of murmann_adc_survey_analyzer using ELDO macromodel
*** This file is parsed to find only the top-level subcircuit
*** Top level subcircuit name is defined with the line below:
*** Design cell name: murmann_adc_survey_analyzer_example

.SUBCKT murmann_adc_survey_analyzer_example IN OUT
    INV0 IN OUT VHI=1 VLO=0 VTHI=0.5 VTLO=0.5 TPD=0.1n
.ENDS
